
module fpga
(
	output 	wire [3:0] pci_exp_txp,
	output 	wire [3:0] pci_exp_txn,

	input 	wire pci_exp_rxp,
	input 	wire pci_exp_rxn,
	input 	wire pcie_refclkin_p,		
	input 	wire pcie_refclkin_n,		
	input 	wire sys_rst_n
		
);


endmodule